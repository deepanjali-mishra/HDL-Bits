// Aim : To assign the constant 0 to the output of a module having 0 inputs and 1 output

module top( output zero ); //Verilog-2001 format
  assign zero = 1'b0;
endmodule
