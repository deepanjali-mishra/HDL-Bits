// Aim: to create a wire  by adding an assign statement to connect in to out

module top_module ( input in, output out );
  assign out = in;
endmodule
