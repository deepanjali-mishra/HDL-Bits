//Aim : To assign logic 1 to output. The module doesn't have any input, and has 1 output

module step_one( output one );
  assign one = 1'b1;
endmodule



