module top_module( input in, output out );
  assign out = ~in; // ~:bitwise not and !: logical not
endmodule
